`include "tb_classes/seq_item.svh"
`include "tb_classes/my_sequence.svh"
`include "tb_classes/driver.svh"
`include "tb_classes/monitor.svh"
`include "tb_classes/sequencer.svh"
`include "tb_classes/agent.svh"
`include "tb_classes/scoreboard.svh"
`include "tb_classes/coverage.svh"
`include "tb_classes/env.svh"
`include "tb_classes/test.svh"